module half_adder(output reg S, output reg C, input wire A, input wire B)



Module full _adder(
input wire [3:0] A
input wire [3:0] B;
input wire[3:0] Cin;
output reg sum;
output reg carry)



half_adder(I1, I2, in1, in2); 
half_adder(sum,I3,I1, cin);

always @